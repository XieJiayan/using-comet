`ifndef AXI_ASSIGN_SVH_
`define AXI_ASSIGN_SVH_



`define AXILITE_ASSIGN(src , dst) 		\
`__AXILITE_TO_AW(assign)



`endif